module register_Q(
input load, //load the register
input rshift, //right shift
input lshift, //left shift
input clk, //clock signal
input right_shift_entry_wire,//signal that enters the register when doing right-shift
input [8:0]qq,//load input bus
input left_shift_entry_wire, //signal that enters the register when doing left-shift
output [8:0]q,//output bus
output [8:0]not_q //inverted output bus
);

wire [1:0]enc;
wire [8:0]d;

encoder4_2 e_inst(.i({lshift, rshift, load, 1'b0}), .o(enc)); //encodes the input signals to an enc bus that goes to the multiplexers as selection signals

genvar i;
generate
	for(i=0;i<=8;i=i+1)
		begin: d_flip_flop
			d_flip_flop d_inst(.d(d[i]), .clk(clk), .q(q[i]), .not_q(not_q[i])); //flip-flops of the register
		end
endgenerate

genvar j; //used 4:2 multiplexers for selecting the input signal for each flip-flop, each of them selects signals in the following order: q[i-1] (when doing left-shift), q[i+1] output (when doing right-shift), load input, q[i] output(memory)
generate
	for(i=0;i<=8;i=i+1)
		begin: mux4_1
			if(i==0)
			mux4_1 mux4_inst0(.i({1'b0, q[i+1], qq[i], q[i]}), .sel(enc), .o(d[i])); //q[0] is used only for multiplication operation, it acts as q[-1] in the booth multiplication algorithm
			else 
			if (i==1)
			mux4_1 mux4_inst1(.i({left_shift_entry_wire, q[i+1], qq[i], q[i]}), .sel(enc), .o(d[i])); //q[1] is used as the least significant bit when doing division, it receives the left shift entry
			else if (i==8)
			mux4_1 mux4_inst2(.i({q[i-1], right_shift_entry_wire, qq[i], q[i]}), .sel(enc), .o(d[i]));
			else
			mux4_1 mux4_inst3(.i({q[i-1], q[i+1], qq[i], q[i]}), .sel(enc), .o(d[i]));//most significant bit
		end
endgenerate

endmodule

module register_Q_tb();

reg load;
reg rshift;
reg lshift;
reg right_shift_entry_wire; 
reg left_shift_entry_wire;
reg clk;
reg [8:0]qq; 
wire [8:0]q; 
wire [8:0]not_q; 

register_Q DUT_REGQ(.load(load), .rshift(rshift), .lshift(lshift), .right_shift_entry_wire(right_shift_entry_wire), .left_shift_entry_wire(left_shift_entry_wire), .clk(clk), .qq(qq), .q(q), .not_q(not_q));

initial begin
clk=1'b0;
repeat (70) #(50) clk=~clk;
end

initial begin
qq=8'b00010111;
load=1;
lshift=0;
rshift=0;
left_shift_entry_wire=0;
right_shift_entry_wire=0;
#100;
qq=8'b01101010;
#100;
load=0;
rshift=1;
#100;
rshift=0;
lshift=1;
left_shift_entry_wire=1;
#400;
lshift=0;
rshift=1;
#400;
rshift=0;
end

endmodule