module mux4_1(input [3:0]i, input [1:0]sel, output o);
	assign o=(i[3]&sel[1]&sel[0]) | (i[2]&sel[1]&~sel[0]) | (i[1]&~sel[1]&sel[0]) | (i[0]&~sel[1]&~sel[0]); 
endmodule